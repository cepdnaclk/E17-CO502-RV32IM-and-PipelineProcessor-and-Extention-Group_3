module alu_int(DATA1, DATA2, SELECT, );

endmodule